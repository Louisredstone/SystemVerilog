module KS_Adder(A,B,Ci,Co,S);
input  [15:0]A;
input  [15:0]B;
input  Ci;
output Co;
output [15:0]S;

wire   [16:0]C;
assign C[0]=Ci;
assign Co=C[16];

wire P_0_0,G_0_0;
wire P_1_1,G_1_1;
wire P_2_2,G_2_2;
wire P_3_3,G_3_3;
wire P_4_4,G_4_4;
wire P_5_5,G_5_5;
wire P_6_6,G_6_6;
wire P_7_7,G_7_7;
wire P_8_8,G_8_8;
wire P_9_9,G_9_9;
wire P_10_10,G_10_10;
wire P_11_11,G_11_11;
wire P_12_12,G_12_12;
wire P_13_13,G_13_13;
wire P_14_14,G_14_14;
wire P_15_15,G_15_15;
wire P_1_0,G_1_0;
wire P_2_1,G_2_1;
wire P_2_0,G_2_0;
wire P_3_2,G_3_2;
wire P_3_0,G_3_0;
wire P_4_3,G_4_3;
wire P_4_1,G_4_1;
wire P_4_0,G_4_0;
wire P_5_4,G_5_4;
wire P_5_2,G_5_2;
wire P_5_0,G_5_0;
wire P_6_5,G_6_5;
wire P_6_3,G_6_3;
wire P_6_0,G_6_0;
wire P_7_6,G_7_6;
wire P_7_4,G_7_4;
wire P_7_0,G_7_0;
wire P_8_7,G_8_7;
wire P_8_5,G_8_5;
wire P_8_1,G_8_1;
wire P_8_0,G_8_0;
wire P_9_8,G_9_8;
wire P_9_6,G_9_6;
wire P_9_2,G_9_2;
wire P_9_0,G_9_0;
wire P_10_9,G_10_9;
wire P_10_7,G_10_7;
wire P_10_3,G_10_3;
wire P_10_0,G_10_0;
wire P_11_10,G_11_10;
wire P_11_8,G_11_8;
wire P_11_4,G_11_4;
wire P_11_0,G_11_0;
wire P_12_11,G_12_11;
wire P_12_9,G_12_9;
wire P_12_5,G_12_5;
wire P_12_0,G_12_0;
wire P_13_12,G_13_12;
wire P_13_10,G_13_10;
wire P_13_6,G_13_6;
wire P_13_0,G_13_0;
wire P_14_13,G_14_13;
wire P_14_11,G_14_11;
wire P_14_7,G_14_7;
wire P_14_0,G_14_0;
wire P_15_14,G_15_14;
wire P_15_12,G_15_12;
wire P_15_8,G_15_8;
wire P_15_0,G_15_0;

assign P_0_0 = A[0] ^ B[0];
assign P_1_1 = A[1] ^ B[1];
assign P_2_2 = A[2] ^ B[2];
assign P_3_3 = A[3] ^ B[3];
assign P_4_4 = A[4] ^ B[4];
assign P_5_5 = A[5] ^ B[5];
assign P_6_6 = A[6] ^ B[6];
assign P_7_7 = A[7] ^ B[7];
assign P_8_8 = A[8] ^ B[8];
assign P_9_9 = A[9] ^ B[9];
assign P_10_10 = A[10] ^ B[10];
assign P_11_11 = A[11] ^ B[11];
assign P_12_12 = A[12] ^ B[12];
assign P_13_13 = A[13] ^ B[13];
assign P_14_14 = A[14] ^ B[14];
assign P_15_15 = A[15] ^ B[15];
assign G_0_0 = A[0] & B[0];
assign G_1_1 = A[1] & B[1];
assign G_2_2 = A[2] & B[2];
assign G_3_3 = A[3] & B[3];
assign G_4_4 = A[4] & B[4];
assign G_5_5 = A[5] & B[5];
assign G_6_6 = A[6] & B[6];
assign G_7_7 = A[7] & B[7];
assign G_8_8 = A[8] & B[8];
assign G_9_9 = A[9] & B[9];
assign G_10_10 = A[10] & B[10];
assign G_11_11 = A[11] & B[11];
assign G_12_12 = A[12] & B[12];
assign G_13_13 = A[13] & B[13];
assign G_14_14 = A[14] & B[14];
assign G_15_15 = A[15] & B[15];

dot dot_1_0(.Pi1(P_1_1),.Gi1(G_1_1),.Pi0(P_0_0),.Gi0(G_0_0),.Po(P_1_0),.Go(G_1_0));
dot dot_2_1(.Pi1(P_2_2),.Gi1(G_2_2),.Pi0(P_1_1),.Gi0(G_1_1),.Po(P_2_1),.Go(G_2_1));
dot dot_2_0(.Pi1(P_2_1),.Gi1(G_2_1),.Pi0(P_0_0),.Gi0(G_0_0),.Po(P_2_0),.Go(G_2_0));
dot dot_3_2(.Pi1(P_3_3),.Gi1(G_3_3),.Pi0(P_2_2),.Gi0(G_2_2),.Po(P_3_2),.Go(G_3_2));
dot dot_3_0(.Pi1(P_3_2),.Gi1(G_3_2),.Pi0(P_1_0),.Gi0(G_1_0),.Po(P_3_0),.Go(G_3_0));
dot dot_4_3(.Pi1(P_4_4),.Gi1(G_4_4),.Pi0(P_3_3),.Gi0(G_3_3),.Po(P_4_3),.Go(G_4_3));
dot dot_4_1(.Pi1(P_4_3),.Gi1(G_4_3),.Pi0(P_2_1),.Gi0(G_2_1),.Po(P_4_1),.Go(G_4_1));
dot dot_4_0(.Pi1(P_4_1),.Gi1(G_4_1),.Pi0(P_0_0),.Gi0(G_0_0),.Po(P_4_0),.Go(G_4_0));
dot dot_5_4(.Pi1(P_5_5),.Gi1(G_5_5),.Pi0(P_4_4),.Gi0(G_4_4),.Po(P_5_4),.Go(G_5_4));
dot dot_5_2(.Pi1(P_5_4),.Gi1(G_5_4),.Pi0(P_3_2),.Gi0(G_3_2),.Po(P_5_2),.Go(G_5_2));
dot dot_5_0(.Pi1(P_5_2),.Gi1(G_5_2),.Pi0(P_1_0),.Gi0(G_1_0),.Po(P_5_0),.Go(G_5_0));
dot dot_6_5(.Pi1(P_6_6),.Gi1(G_6_6),.Pi0(P_5_5),.Gi0(G_5_5),.Po(P_6_5),.Go(G_6_5));
dot dot_6_3(.Pi1(P_6_5),.Gi1(G_6_5),.Pi0(P_4_3),.Gi0(G_4_3),.Po(P_6_3),.Go(G_6_3));
dot dot_6_0(.Pi1(P_6_3),.Gi1(G_6_3),.Pi0(P_2_0),.Gi0(G_2_0),.Po(P_6_0),.Go(G_6_0));
dot dot_7_6(.Pi1(P_7_7),.Gi1(G_7_7),.Pi0(P_6_6),.Gi0(G_6_6),.Po(P_7_6),.Go(G_7_6));
dot dot_7_4(.Pi1(P_7_6),.Gi1(G_7_6),.Pi0(P_5_4),.Gi0(G_5_4),.Po(P_7_4),.Go(G_7_4));
dot dot_7_0(.Pi1(P_7_4),.Gi1(G_7_4),.Pi0(P_3_0),.Gi0(G_3_0),.Po(P_7_0),.Go(G_7_0));
dot dot_8_7(.Pi1(P_8_8),.Gi1(G_8_8),.Pi0(P_7_7),.Gi0(G_7_7),.Po(P_8_7),.Go(G_8_7));
dot dot_8_5(.Pi1(P_8_7),.Gi1(G_8_7),.Pi0(P_6_5),.Gi0(G_6_5),.Po(P_8_5),.Go(G_8_5));
dot dot_8_1(.Pi1(P_8_5),.Gi1(G_8_5),.Pi0(P_4_1),.Gi0(G_4_1),.Po(P_8_1),.Go(G_8_1));
dot dot_8_0(.Pi1(P_8_1),.Gi1(G_8_1),.Pi0(P_0_0),.Gi0(G_0_0),.Po(P_8_0),.Go(G_8_0));
dot dot_9_8(.Pi1(P_9_9),.Gi1(G_9_9),.Pi0(P_8_8),.Gi0(G_8_8),.Po(P_9_8),.Go(G_9_8));
dot dot_9_6(.Pi1(P_9_8),.Gi1(G_9_8),.Pi0(P_7_6),.Gi0(G_7_6),.Po(P_9_6),.Go(G_9_6));
dot dot_9_2(.Pi1(P_9_6),.Gi1(G_9_6),.Pi0(P_5_2),.Gi0(G_5_2),.Po(P_9_2),.Go(G_9_2));
dot dot_9_0(.Pi1(P_9_2),.Gi1(G_9_2),.Pi0(P_1_0),.Gi0(G_1_0),.Po(P_9_0),.Go(G_9_0));
dot dot_10_9(.Pi1(P_10_10),.Gi1(G_10_10),.Pi0(P_9_9),.Gi0(G_9_9),.Po(P_10_9),.Go(G_10_9));
dot dot_10_7(.Pi1(P_10_9),.Gi1(G_10_9),.Pi0(P_8_7),.Gi0(G_8_7),.Po(P_10_7),.Go(G_10_7));
dot dot_10_3(.Pi1(P_10_7),.Gi1(G_10_7),.Pi0(P_6_3),.Gi0(G_6_3),.Po(P_10_3),.Go(G_10_3));
dot dot_10_0(.Pi1(P_10_3),.Gi1(G_10_3),.Pi0(P_2_0),.Gi0(G_2_0),.Po(P_10_0),.Go(G_10_0));
dot dot_11_10(.Pi1(P_11_11),.Gi1(G_11_11),.Pi0(P_10_10),.Gi0(G_10_10),.Po(P_11_10),.Go(G_11_10));
dot dot_11_8(.Pi1(P_11_10),.Gi1(G_11_10),.Pi0(P_9_8),.Gi0(G_9_8),.Po(P_11_8),.Go(G_11_8));
dot dot_11_4(.Pi1(P_11_8),.Gi1(G_11_8),.Pi0(P_7_4),.Gi0(G_7_4),.Po(P_11_4),.Go(G_11_4));
dot dot_11_0(.Pi1(P_11_4),.Gi1(G_11_4),.Pi0(P_3_0),.Gi0(G_3_0),.Po(P_11_0),.Go(G_11_0));
dot dot_12_11(.Pi1(P_12_12),.Gi1(G_12_12),.Pi0(P_11_11),.Gi0(G_11_11),.Po(P_12_11),.Go(G_12_11));
dot dot_12_9(.Pi1(P_12_11),.Gi1(G_12_11),.Pi0(P_10_9),.Gi0(G_10_9),.Po(P_12_9),.Go(G_12_9));
dot dot_12_5(.Pi1(P_12_9),.Gi1(G_12_9),.Pi0(P_8_5),.Gi0(G_8_5),.Po(P_12_5),.Go(G_12_5));
dot dot_12_0(.Pi1(P_12_5),.Gi1(G_12_5),.Pi0(P_4_0),.Gi0(G_4_0),.Po(P_12_0),.Go(G_12_0));
dot dot_13_12(.Pi1(P_13_13),.Gi1(G_13_13),.Pi0(P_12_12),.Gi0(G_12_12),.Po(P_13_12),.Go(G_13_12));
dot dot_13_10(.Pi1(P_13_12),.Gi1(G_13_12),.Pi0(P_11_10),.Gi0(G_11_10),.Po(P_13_10),.Go(G_13_10));
dot dot_13_6(.Pi1(P_13_10),.Gi1(G_13_10),.Pi0(P_9_6),.Gi0(G_9_6),.Po(P_13_6),.Go(G_13_6));
dot dot_13_0(.Pi1(P_13_6),.Gi1(G_13_6),.Pi0(P_5_0),.Gi0(G_5_0),.Po(P_13_0),.Go(G_13_0));
dot dot_14_13(.Pi1(P_14_14),.Gi1(G_14_14),.Pi0(P_13_13),.Gi0(G_13_13),.Po(P_14_13),.Go(G_14_13));
dot dot_14_11(.Pi1(P_14_13),.Gi1(G_14_13),.Pi0(P_12_11),.Gi0(G_12_11),.Po(P_14_11),.Go(G_14_11));
dot dot_14_7(.Pi1(P_14_11),.Gi1(G_14_11),.Pi0(P_10_7),.Gi0(G_10_7),.Po(P_14_7),.Go(G_14_7));
dot dot_14_0(.Pi1(P_14_7),.Gi1(G_14_7),.Pi0(P_6_0),.Gi0(G_6_0),.Po(P_14_0),.Go(G_14_0));
dot dot_15_14(.Pi1(P_15_15),.Gi1(G_15_15),.Pi0(P_14_14),.Gi0(G_14_14),.Po(P_15_14),.Go(G_15_14));
dot dot_15_12(.Pi1(P_15_14),.Gi1(G_15_14),.Pi0(P_13_12),.Gi0(G_13_12),.Po(P_15_12),.Go(G_15_12));
dot dot_15_8(.Pi1(P_15_12),.Gi1(G_15_12),.Pi0(P_11_8),.Gi0(G_11_8),.Po(P_15_8),.Go(G_15_8));
dot dot_15_0(.Pi1(P_15_8),.Gi1(G_15_8),.Pi0(P_7_0),.Gi0(G_7_0),.Po(P_15_0),.Go(G_15_0));

assign C[1] = G_0_0 | (P_0_0 & C[0]);
assign C[2] = G_1_0 | (P_1_0 & C[0]);
assign C[3] = G_2_0 | (P_2_0 & C[0]);
assign C[4] = G_3_0 | (P_3_0 & C[0]);
assign C[5] = G_4_0 | (P_4_0 & C[0]);
assign C[6] = G_5_0 | (P_5_0 & C[0]);
assign C[7] = G_6_0 | (P_6_0 & C[0]);
assign C[8] = G_7_0 | (P_7_0 & C[0]);
assign C[9] = G_8_0 | (P_8_0 & C[0]);
assign C[10] = G_9_0 | (P_9_0 & C[0]);
assign C[11] = G_10_0 | (P_10_0 & C[0]);
assign C[12] = G_11_0 | (P_11_0 & C[0]);
assign C[13] = G_12_0 | (P_12_0 & C[0]);
assign C[14] = G_13_0 | (P_13_0 & C[0]);
assign C[15] = G_14_0 | (P_14_0 & C[0]);
assign C[16] = G_15_0 | (P_15_0 & C[0]);

assign S[0] = P_0_0 ^ C[0];
assign S[1] = P_1_1 ^ C[1];
assign S[2] = P_2_2 ^ C[2];
assign S[3] = P_3_3 ^ C[3];
assign S[4] = P_4_4 ^ C[4];
assign S[5] = P_5_5 ^ C[5];
assign S[6] = P_6_6 ^ C[6];
assign S[7] = P_7_7 ^ C[7];
assign S[8] = P_8_8 ^ C[8];
assign S[9] = P_9_9 ^ C[9];
assign S[10] = P_10_10 ^ C[10];
assign S[11] = P_11_11 ^ C[11];
assign S[12] = P_12_12 ^ C[12];
assign S[13] = P_13_13 ^ C[13];
assign S[14] = P_14_14 ^ C[14];
assign S[15] = P_15_15 ^ C[15];

endmodule

module dot(Pi1,Gi1,Pi0,Gi0,Po,Go);
//P"i:j" = P"i:m" & P"m-1:j"
//G"i:j" = G"i:m" | P"i:m" & G"m-i:j"
//Pi0: P"m-1:j"
//Gi0: G"m-1:j"
//Pi1: P"i:m"
//Gi1: G"i:m"
//Po:  P"i:j"
//Go:  G"i:j"
input  Pi0,Gi0,Pi1,Gi1;
output Po,Go;

assign Po = Pi1 & Pi0;
assign Go = Gi1 | (Pi1 & Gi0);
endmodule
